module pipeemreg (ewreg,em2reg,ewmem,ealu,eb,ern,clock,resetn,
							mwreg,mm2reg,mwmem,malu,mb,mrn); // EXE/MEM流水线寄存器

//EXE/MEM流水线寄存器模块，起承接EXE阶段和MEM阶段的流水任务。 
//在 clock 上升沿时，将 EXE 阶段需传递给MEM阶段的信息，锁存在EXE/MEM 
//流水线寄存器中，并呈现在MEM阶段。 

input           ewreg, em2reg, ewmem, clock, resetn;
input [31:0]    ealu, eb; 
input [4:0]     ern;

output          mwreg, mm2reg, mwmem;
output [31:0]   malu, mb; 
output [4:0]    mrn;


reg          mwreg, mm2reg, mwmem;
reg [31:0]   malu, mb; 
reg [4:0]    mrn;
always @ (negedge resetn or posedge clock)
      if (resetn == 0) 
         begin
            malu       <= 32'b0;
            mb         <= 32'b0;
            mrn        <=  4'b0;
            mwreg      <=  1'b0;
            mm2reg     <=  1'b0;
            mwmem      <=  1'b0;
         end 
      else
         begin 
            malu       <= ealu;
            mb         <= eb;
            mrn        <= ern;
            mwreg      <= ewreg;
            mm2reg     <= em2reg;
            mwmem      <= ewmem;
         end
endmodule
